// DE2_115_SOPC.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		input  wire        vid_clk_to_the_alt_vip_itc_0,             //         alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] vid_data_from_the_alt_vip_itc_0,          //                                    .vid_data
		output wire        underflow_from_the_alt_vip_itc_0,         //                                    .underflow
		output wire        vid_datavalid_from_the_alt_vip_itc_0,     //                                    .vid_datavalid
		output wire        vid_v_sync_from_the_alt_vip_itc_0,        //                                    .vid_v_sync
		output wire        vid_h_sync_from_the_alt_vip_itc_0,        //                                    .vid_h_sync
		output wire        vid_f_from_the_alt_vip_itc_0,             //                                    .vid_f
		output wire        vid_h_from_the_alt_vip_itc_0,             //                                    .vid_h
		output wire        vid_v_from_the_alt_vip_itc_0,             //                                    .vid_v
		input  wire        altpll_0_areset_conduit_export,           //             altpll_0_areset_conduit.export
		output wire        altpll_0_c1_out,                          //                         altpll_0_c1.clk
		output wire        locked_from_the_altpll_0,                 //             altpll_0_locked_conduit.export
		output wire        phasedone_from_the_altpll_0,              //          altpll_0_phasedone_conduit.export
		output wire        altpll_audio_locked_conduit_export,       //         altpll_audio_locked_conduit.export
		output wire        altpll_audio_phasedone_conduit_export,    //      altpll_audio_phasedone_conduit.export
		output wire        audio_conduit_end_XCK,                    //                   audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                 //                                    .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                 //                                    .ADCLRC
		output wire        audio_conduit_end_DACDAT,                 //                                    .DACDAT
		input  wire        audio_conduit_end_DACLRC,                 //                                    .DACLRC
		input  wire        audio_conduit_end_BCLK,                   //                                    .BCLK
		input  wire        clk_50,                                   //                       clk_50_clk_in.clk
		input  wire        reset_n,                                  //                 clk_50_clk_in_reset.reset_n
		output wire        dclk_from_the_epcs_flash_controller,      //      epcs_flash_controller_external.dclk
		output wire        sce_from_the_epcs_flash_controller,       //                                    .sce
		output wire        sdo_from_the_epcs_flash_controller,       //                                    .sdo
		input  wire        data0_to_the_epcs_flash_controller,       //                                    .data0
		inout  wire        i2c_opencores_0_export_scl_pad_io,        //              i2c_opencores_0_export.scl_pad_io
		inout  wire        i2c_opencores_0_export_sda_pad_io,        //                                    .sda_pad_io
		output wire        i2c_scl_external_connection_export,       //         i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,       //         i2c_sda_external_connection.export
		input  wire [3:0]  in_port_to_the_key,                       //             key_external_connection.export
		output wire        LCD_RS_from_the_lcd,                      //                        lcd_external.RS
		output wire        LCD_RW_from_the_lcd,                      //                                    .RW
		inout  wire [7:0]  LCD_data_to_and_from_the_lcd,             //                                    .data
		output wire        LCD_E_from_the_lcd,                       //                                    .E
		input  wire        lcd_touch_int_external_connection_export, //   lcd_touch_int_external_connection.export
		output wire [26:0] out_port_from_the_led,                    //             led_external_connection.export
		output wire        sd_clk_external_connection_export,        //          sd_clk_external_connection.export
		inout  wire        sd_cmd_external_connection_export,        //          sd_cmd_external_connection.export
		inout  wire [3:0]  sd_dat_external_connection_export,        //          sd_dat_external_connection.export
		input  wire        sd_wp_n_external_connection_export,       //         sd_wp_n_external_connection.export
		output wire [12:0] zs_addr_from_the_sdram,                   //                          sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                     //                                    .ba
		output wire        zs_cas_n_from_the_sdram,                  //                                    .cas_n
		output wire        zs_cke_from_the_sdram,                    //                                    .cke
		output wire        zs_cs_n_from_the_sdram,                   //                                    .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram,              //                                    .dq
		output wire [3:0]  zs_dqm_from_the_sdram,                    //                                    .dqm
		output wire        zs_ras_n_from_the_sdram,                  //                                    .ras_n
		output wire        zs_we_n_from_the_sdram,                   //                                    .we_n
		inout  wire [15:0] SRAM_DQ_to_and_from_the_sram,             //                    sram_conduit_end.DQ
		output wire [19:0] SRAM_ADDR_from_the_sram,                  //                                    .ADDR
		output wire        SRAM_UB_n_from_the_sram,                  //                                    .UB_n
		output wire        SRAM_LB_n_from_the_sram,                  //                                    .LB_n
		output wire        SRAM_WE_n_from_the_sram,                  //                                    .WE_n
		output wire        SRAM_CE_n_from_the_sram,                  //                                    .CE_n
		output wire        SRAM_OE_n_from_the_sram,                  //                                    .OE_n
		input  wire [17:0] in_port_to_the_sw,                        //              sw_external_connection.export
		inout  wire [7:0]  data_to_and_from_the_cfi_flash,           // tri_state_bridge_flash_bridge_0_out.data_to_and_from_the_cfi_flash
		output wire [22:0] address_to_the_cfi_flash,                 //                                    .address_to_the_cfi_flash
		output wire [0:0]  write_n_to_the_cfi_flash,                 //                                    .write_n_to_the_cfi_flash
		output wire [0:0]  select_n_to_the_cfi_flash,                //                                    .select_n_to_the_cfi_flash
		output wire [0:0]  read_n_to_the_cfi_flash                   //                                    .read_n_to_the_cfi_flash
	);

	wire         alt_vip_vfr_0_avalon_streaming_source_valid;                                 // alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	wire  [23:0] alt_vip_vfr_0_avalon_streaming_source_data;                                  // alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	wire         alt_vip_vfr_0_avalon_streaming_source_ready;                                 // alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	wire         alt_vip_vfr_0_avalon_streaming_source_startofpacket;                         // alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire         alt_vip_vfr_0_avalon_streaming_source_endofpacket;                           // alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire         altpll_0_c0_clk;                                                             // altpll_0:c0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_0:clock, alt_vip_vfr_0:master_clock, cfi_flash:clk_clk, clock_crossing_io:s0_clk, cpu:clk, epcs_flash_controller:clk, i2c_scl:clk, i2c_sda:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, jtag_uart:clk, key:clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, rst_controller:clk, rst_controller_006:clk, sd_clk:clk, sd_cmd:clk, sd_dat:clk, sd_wp_n:clk, sdram:clk, sram:clk, tri_state_bridge_flash_bridge_0:clk, tri_state_bridge_flash_pinSharer_0:clk_clk]
	wire         altpll_audio_c0_clk;                                                         // altpll_audio:c0 -> [audio:avs_s1_clk, mm_interconnect_0:altpll_audio_c0_clk, rst_controller_003:clk]
	wire         altpll_0_c2_clk;                                                             // altpll_0:c2 -> [clock_crossing_io:m0_clk, irq_synchronizer_001:receiver_clk, lcd:clk, led:clk, mm_interconnect_1:altpll_0_c2_clk, rst_controller_004:clk, sw:clk, sysid:clock, timer:clk]
	wire         altpll_0_c3_clk;                                                             // altpll_0:c3 -> [i2c_opencores_0:wb_clk_i, irq_synchronizer:receiver_clk, irq_synchronizer_002:receiver_clk, lcd_touch_int:clk, mm_interconnect_0:altpll_0_c3_clk, rst_controller_005:clk]
	wire         tri_state_bridge_flash_pinsharer_0_tcm_request;                              // tri_state_bridge_flash_pinSharer_0:request -> tri_state_bridge_flash_bridge_0:request
	wire   [7:0] tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_in;    // tri_state_bridge_flash_bridge_0:tcs_data_to_and_from_the_cfi_flash_in -> tri_state_bridge_flash_pinSharer_0:data_to_and_from_the_cfi_flash_in
	wire   [0:0] tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out;          // tri_state_bridge_flash_pinSharer_0:read_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_read_n_to_the_cfi_flash
	wire  [22:0] tri_state_bridge_flash_pinsharer_0_tcm_address_to_the_cfi_flash_out;         // tri_state_bridge_flash_pinSharer_0:address_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_address_to_the_cfi_flash
	wire   [7:0] tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_out;   // tri_state_bridge_flash_pinSharer_0:data_to_and_from_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_data_to_and_from_the_cfi_flash
	wire   [0:0] tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out;         // tri_state_bridge_flash_pinSharer_0:write_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_write_n_to_the_cfi_flash
	wire         tri_state_bridge_flash_pinsharer_0_tcm_grant;                                // tri_state_bridge_flash_bridge_0:grant -> tri_state_bridge_flash_pinSharer_0:grant
	wire         tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_outen; // tri_state_bridge_flash_pinSharer_0:data_to_and_from_the_cfi_flash_outen -> tri_state_bridge_flash_bridge_0:tcs_data_to_and_from_the_cfi_flash_outen
	wire   [0:0] tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out;        // tri_state_bridge_flash_pinSharer_0:select_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_select_n_to_the_cfi_flash
	wire         cfi_flash_tcm_data_outen;                                                    // cfi_flash:tcm_data_outen -> tri_state_bridge_flash_pinSharer_0:tcs0_data_outen
	wire         cfi_flash_tcm_request;                                                       // cfi_flash:tcm_request -> tri_state_bridge_flash_pinSharer_0:tcs0_request
	wire         cfi_flash_tcm_write_n_out;                                                   // cfi_flash:tcm_write_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_write_n_out
	wire         cfi_flash_tcm_read_n_out;                                                    // cfi_flash:tcm_read_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_read_n_out
	wire         cfi_flash_tcm_grant;                                                         // tri_state_bridge_flash_pinSharer_0:tcs0_grant -> cfi_flash:tcm_grant
	wire         cfi_flash_tcm_chipselect_n_out;                                              // cfi_flash:tcm_chipselect_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_chipselect_n_out
	wire  [22:0] cfi_flash_tcm_address_out;                                                   // cfi_flash:tcm_address_out -> tri_state_bridge_flash_pinSharer_0:tcs0_address_out
	wire   [7:0] cfi_flash_tcm_data_out;                                                      // cfi_flash:tcm_data_out -> tri_state_bridge_flash_pinSharer_0:tcs0_data_out
	wire   [7:0] cfi_flash_tcm_data_in;                                                       // tri_state_bridge_flash_pinSharer_0:tcs0_data_in -> cfi_flash:tcm_data_in
	wire  [31:0] alt_vip_vfr_0_avalon_master_readdata;                                        // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire         alt_vip_vfr_0_avalon_master_waitrequest;                                     // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire  [31:0] alt_vip_vfr_0_avalon_master_address;                                         // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire         alt_vip_vfr_0_avalon_master_read;                                            // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire         alt_vip_vfr_0_avalon_master_readdatavalid;                                   // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire   [5:0] alt_vip_vfr_0_avalon_master_burstcount;                                      // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire  [31:0] cpu_data_master_readdata;                                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                               // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_sdram_s1_chipselect;                                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_sram_avalon_slave_chipselect;                              // mm_interconnect_0:sram_avalon_slave_chipselect -> sram:s_chipselect_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_readdata;                                // sram:s_readdata -> mm_interconnect_0:sram_avalon_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_slave_address;                                 // mm_interconnect_0:sram_avalon_slave_address -> sram:s_address
	wire         mm_interconnect_0_sram_avalon_slave_read;                                    // mm_interconnect_0:sram_avalon_slave_read -> sram:s_read_n
	wire   [1:0] mm_interconnect_0_sram_avalon_slave_byteenable;                              // mm_interconnect_0:sram_avalon_slave_byteenable -> sram:s_byteenable_n
	wire         mm_interconnect_0_sram_avalon_slave_write;                                   // mm_interconnect_0:sram_avalon_slave_write -> sram:s_write_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_writedata;                               // mm_interconnect_0:sram_avalon_slave_writedata -> sram:s_writedata
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata;                       // alt_vip_vfr_0:slave_readdata -> mm_interconnect_0:alt_vip_vfr_0_avalon_slave_readdata
	wire   [4:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address;                        // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read;                           // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write;                          // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata;                      // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_readdata;                               // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_audio_avalon_slave_address;                                // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire         mm_interconnect_0_audio_avalon_slave_read;                                   // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire         mm_interconnect_0_audio_avalon_slave_write;                                  // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_writedata;                              // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect;                 // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata;                   // i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest;                // i2c_opencores_0:wb_ack_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address;                    // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write;                      // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata;                  // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect;        // mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata;          // epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_address;           // mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;              // mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> epcs_flash_controller:read_n
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;             // mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> epcs_flash_controller:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata;         // mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                               // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                                   // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                                  // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                              // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_readdata;                           // altpll_audio:readdata -> mm_interconnect_0:altpll_audio_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_audio_pll_slave_address;                            // mm_interconnect_0:altpll_audio_pll_slave_address -> altpll_audio:address
	wire         mm_interconnect_0_altpll_audio_pll_slave_read;                               // mm_interconnect_0:altpll_audio_pll_slave_read -> altpll_audio:read
	wire         mm_interconnect_0_altpll_audio_pll_slave_write;                              // mm_interconnect_0:altpll_audio_pll_slave_write -> altpll_audio:write
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_writedata;                          // mm_interconnect_0:altpll_audio_pll_slave_writedata -> altpll_audio:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                             // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                          // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                          // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire   [8:0] mm_interconnect_0_clock_crossing_io_s0_address;                              // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                                 // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                           // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                        // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                                // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                            // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                           // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_lcd_touch_int_s1_chipselect;                               // mm_interconnect_0:lcd_touch_int_s1_chipselect -> lcd_touch_int:chipselect
	wire  [31:0] mm_interconnect_0_lcd_touch_int_s1_readdata;                                 // lcd_touch_int:readdata -> mm_interconnect_0:lcd_touch_int_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_touch_int_s1_address;                                  // mm_interconnect_0:lcd_touch_int_s1_address -> lcd_touch_int:address
	wire         mm_interconnect_0_lcd_touch_int_s1_write;                                    // mm_interconnect_0:lcd_touch_int_s1_write -> lcd_touch_int:write_n
	wire  [31:0] mm_interconnect_0_lcd_touch_int_s1_writedata;                                // mm_interconnect_0:lcd_touch_int_s1_writedata -> lcd_touch_int:writedata
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_readdata;                                    // cfi_flash:uas_readdata -> mm_interconnect_0:cfi_flash_uas_readdata
	wire         mm_interconnect_0_cfi_flash_uas_waitrequest;                                 // cfi_flash:uas_waitrequest -> mm_interconnect_0:cfi_flash_uas_waitrequest
	wire         mm_interconnect_0_cfi_flash_uas_debugaccess;                                 // mm_interconnect_0:cfi_flash_uas_debugaccess -> cfi_flash:uas_debugaccess
	wire  [22:0] mm_interconnect_0_cfi_flash_uas_address;                                     // mm_interconnect_0:cfi_flash_uas_address -> cfi_flash:uas_address
	wire         mm_interconnect_0_cfi_flash_uas_read;                                        // mm_interconnect_0:cfi_flash_uas_read -> cfi_flash:uas_read
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_byteenable;                                  // mm_interconnect_0:cfi_flash_uas_byteenable -> cfi_flash:uas_byteenable
	wire         mm_interconnect_0_cfi_flash_uas_readdatavalid;                               // cfi_flash:uas_readdatavalid -> mm_interconnect_0:cfi_flash_uas_readdatavalid
	wire         mm_interconnect_0_cfi_flash_uas_lock;                                        // mm_interconnect_0:cfi_flash_uas_lock -> cfi_flash:uas_lock
	wire         mm_interconnect_0_cfi_flash_uas_write;                                       // mm_interconnect_0:cfi_flash_uas_write -> cfi_flash:uas_write
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_writedata;                                   // mm_interconnect_0:cfi_flash_uas_writedata -> cfi_flash:uas_writedata
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_burstcount;                                  // mm_interconnect_0:cfi_flash_uas_burstcount -> cfi_flash:uas_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                            // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                                               // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                            // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [8:0] clock_crossing_io_m0_address;                                                // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                                   // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                                             // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                          // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                                              // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                                  // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                                             // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;                                // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;                                 // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_read;                                    // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;                           // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_1_lcd_control_slave_write;                                   // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;                               // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                              // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                               // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_timer_s1_chipselect;                                       // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                         // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                          // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                                            // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                        // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_1_led_s1_chipselect;                                         // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                           // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                            // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                                              // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                          // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                            // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                             // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_key_s1_chipselect;                                         // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                           // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                            // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                                              // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                          // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_sd_clk_s1_chipselect;                                      // mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	wire  [31:0] mm_interconnect_1_sd_clk_s1_readdata;                                        // sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_clk_s1_address;                                         // mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	wire         mm_interconnect_1_sd_clk_s1_write;                                           // mm_interconnect_1:sd_clk_s1_write -> sd_clk:write_n
	wire  [31:0] mm_interconnect_1_sd_clk_s1_writedata;                                       // mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	wire         mm_interconnect_1_sd_cmd_s1_chipselect;                                      // mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_readdata;                                        // sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_cmd_s1_address;                                         // mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	wire         mm_interconnect_1_sd_cmd_s1_write;                                           // mm_interconnect_1:sd_cmd_s1_write -> sd_cmd:write_n
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_writedata;                                       // mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	wire         mm_interconnect_1_sd_dat_s1_chipselect;                                      // mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	wire  [31:0] mm_interconnect_1_sd_dat_s1_readdata;                                        // sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_dat_s1_address;                                         // mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	wire         mm_interconnect_1_sd_dat_s1_write;                                           // mm_interconnect_1:sd_dat_s1_write -> sd_dat:write_n
	wire  [31:0] mm_interconnect_1_sd_dat_s1_writedata;                                       // mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	wire  [31:0] mm_interconnect_1_sd_wp_n_s1_readdata;                                       // sd_wp_n:readdata -> mm_interconnect_1:sd_wp_n_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_wp_n_s1_address;                                        // mm_interconnect_1:sd_wp_n_s1_address -> sd_wp_n:address
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                                     // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                                       // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                                        // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_write;                                          // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                                      // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                                     // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                                       // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                                        // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_write;                                          // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                                      // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire         irq_mapper_receiver0_irq;                                                    // alt_vip_vfr_0:slave_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver2_irq;                                                    // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver4_irq;                                                    // key:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                    // epcs_flash_controller:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_irq_irq;                                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver1_irq;                                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                               // i2c_opencores_0:wb_inta_o -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                           // timer:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver6_irq;                                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                           // lcd_touch_int:irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_0:master_reset, alt_vip_vfr_0:reset, cfi_flash:reset_reset, clock_crossing_io:s0_reset, cpu:reset_n, epcs_flash_controller:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, key:reset_n, mm_interconnect_0:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_1:key_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sram:reset_n, tri_state_bridge_flash_bridge_0:reset, tri_state_bridge_flash_pinSharer_0:reset_reset]
	wire         rst_controller_reset_out_reset_req;                                          // rst_controller:reset_req -> [cpu:reset_req, epcs_flash_controller:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                               // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_004:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                          // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                          // rst_controller_002:reset_out -> [altpll_audio:reset, mm_interconnect_0:altpll_audio_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                          // rst_controller_003:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_clock_sink_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                                          // rst_controller_004:reset_out -> [clock_crossing_io:m0_reset, irq_synchronizer_001:receiver_reset, lcd:reset_n, led:reset_n, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, sw:reset_n, sysid:reset_n, timer:reset_n]
	wire         rst_controller_005_reset_out_reset;                                          // rst_controller_005:reset_out -> [i2c_opencores_0:wb_rst_i, irq_synchronizer:receiver_reset, irq_synchronizer_002:receiver_reset, lcd_touch_int:reset_n, mm_interconnect_0:i2c_opencores_0_clock_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_006_reset_out_reset;                                          // rst_controller_006:reset_out -> [i2c_scl:reset_n, i2c_sda:reset_n, mm_interconnect_1:sd_clk_reset_reset_bridge_in_reset_reset, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, sd_wp_n:reset_n]

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (800),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (800),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (799),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (30),
		.H_FRONT_PORCH                 (210),
		.H_BACK_PORCH                  (16),
		.V_SYNC_LENGTH                 (13),
		.V_FRONT_PORCH                 (22),
		.V_BACK_PORCH                  (10),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (altpll_0_c0_clk),                                     //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),                      // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (vid_clk_to_the_alt_vip_itc_0),                        //    clocked_video.export
		.vid_data      (vid_data_from_the_alt_vip_itc_0),                     //                 .export
		.underflow     (underflow_from_the_alt_vip_itc_0),                    //                 .export
		.vid_datavalid (vid_datavalid_from_the_alt_vip_itc_0),                //                 .export
		.vid_v_sync    (vid_v_sync_from_the_alt_vip_itc_0),                   //                 .export
		.vid_h_sync    (vid_h_sync_from_the_alt_vip_itc_0),                   //                 .export
		.vid_f         (vid_f_from_the_alt_vip_itc_0),                        //                 .export
		.vid_h         (vid_h_from_the_alt_vip_itc_0),                        //                 .export
		.vid_v         (vid_v_from_the_alt_vip_itc_0)                         //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (800),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (0)
	) alt_vip_vfr_0 (
		.clock                (altpll_0_c0_clk),                                        //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (altpll_0_c0_clk),                                        //            clock_master.clk
		.master_reset         (rst_controller_reset_out_reset),                         //      clock_master_reset.reset
		.slave_address        (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (irq_mapper_receiver0_irq),                               //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	DE2_115_SOPC_altpll_0 altpll_0 (
		.clk       (clk_50),                                         //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                //                    c0.clk
		.c1        (altpll_0_c1_out),                                //                    c1.clk
		.c2        (altpll_0_c2_clk),                                //                    c2.clk
		.c3        (altpll_0_c3_clk),                                //                    c3.clk
		.areset    (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked    (locked_from_the_altpll_0),                       //        locked_conduit.export
		.phasedone (phasedone_from_the_altpll_0)                     //     phasedone_conduit.export
	);

	DE2_115_SOPC_altpll_audio altpll_audio (
		.clk       (clk_50),                                             //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),                 // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_audio_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_audio_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_audio_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_audio_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_audio_pll_slave_writedata), //                      .writedata
		.c0        (altpll_audio_c0_clk),                                //                    c0.clk
		.areset    (),                                                   //        areset_conduit.export
		.locked    (altpll_audio_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_audio_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	AUDIO_IF audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (altpll_audio_c0_clk),                            //       clock_sink.clk
		.avs_s1_reset         (rst_controller_003_reset_out_reset),             // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	DE2_115_SOPC_cfi_flash #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash (
		.clk_clk              (altpll_0_c0_clk),                               //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                // reset.reset
		.uas_address          (mm_interconnect_0_cfi_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_cfi_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_cfi_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_cfi_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_cfi_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_cfi_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_cfi_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_cfi_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_cfi_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_cfi_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_cfi_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (cfi_flash_tcm_request),                         //      .request
		.tcm_grant            (cfi_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (cfi_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (cfi_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (cfi_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (cfi_flash_tcm_data_in)                          //      .data_in
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_0_c2_clk),                                      //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                                      //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                 (altpll_0_c0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DE2_115_SOPC_epcs_flash_controller epcs_flash_controller (
		.clk           (altpll_0_c0_clk),                                                      //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                      //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                                   //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                                     //                  .dataavailable
		.endofpacket   (),                                                                     //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                                     //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver5_irq),                                             //               irq.irq
		.dclk          (dclk_from_the_epcs_flash_controller),                                  //          external.export
		.sce           (sce_from_the_epcs_flash_controller),                                   //                  .export
		.sdo           (sdo_from_the_epcs_flash_controller),                                   //                  .export
		.data0         (data0_to_the_epcs_flash_controller)                                    //                  .export
	);

	i2c_opencores i2c_opencores_0 (
		.wb_clk_i   (altpll_0_c3_clk),                                              //            clock.clk
		.wb_rst_i   (rst_controller_005_reset_out_reset),                           //      clock_reset.reset
		.scl_pad_io (i2c_opencores_0_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_0_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_receiver_irq)                                 // interrupt_sender.irq
	);

	DE2_115_SOPC_i2c_scl i2c_scl (
		.clk        (altpll_0_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_sda i2c_sda (
		.clk        (altpll_0_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_0_c0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	DE2_115_SOPC_key key (
		.clk        (altpll_0_c0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_mapper_receiver4_irq)             //                 irq.irq
	);

	DE2_115_SOPC_lcd lcd (
		.reset_n       (~rst_controller_004_reset_out_reset),               //         reset.reset_n
		.clk           (altpll_0_c2_clk),                                   //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (LCD_RS_from_the_lcd),                               //      external.export
		.LCD_RW        (LCD_RW_from_the_lcd),                               //              .export
		.LCD_data      (LCD_data_to_and_from_the_lcd),                      //              .export
		.LCD_E         (LCD_E_from_the_lcd)                                 //              .export
	);

	DE2_115_SOPC_lcd_touch_int lcd_touch_int (
		.clk        (altpll_0_c3_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_lcd_touch_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_touch_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_touch_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_touch_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_touch_int_s1_readdata),   //                    .readdata
		.in_port    (lcd_touch_int_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)              //                 irq.irq
	);

	DE2_115_SOPC_led led (
		.clk        (altpll_0_c2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led)                // external_connection.export
	);

	DE2_115_SOPC_i2c_scl sd_clk (
		.clk        (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_sda sd_cmd (
		.clk        (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sd_dat sd_dat (
		.clk        (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sd_wp_n sd_wp_n (
		.clk      (altpll_0_c0_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_006_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_1_sd_wp_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sd_wp_n_s1_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)     // external_connection.export
	);

	DE2_115_SOPC_sdram sdram (
		.clk            (altpll_0_c0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (altpll_0_c0_clk),                                 //       clock_reset.clk
		.reset_n        (~rst_controller_reset_out_reset),                 // clock_reset_reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_sram_avalon_slave_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~mm_interconnect_0_sram_avalon_slave_write),      //                  .write_n
		.s_address      (mm_interconnect_0_sram_avalon_slave_address),     //                  .address
		.s_read_n       (~mm_interconnect_0_sram_avalon_slave_read),       //                  .read_n
		.s_writedata    (mm_interconnect_0_sram_avalon_slave_writedata),   //                  .writedata
		.s_readdata     (mm_interconnect_0_sram_avalon_slave_readdata),    //                  .readdata
		.s_byteenable_n (~mm_interconnect_0_sram_avalon_slave_byteenable), //                  .byteenable_n
		.SRAM_DQ        (SRAM_DQ_to_and_from_the_sram),                    //       conduit_end.export
		.SRAM_ADDR      (SRAM_ADDR_from_the_sram),                         //                  .export
		.SRAM_UB_n      (SRAM_UB_n_from_the_sram),                         //                  .export
		.SRAM_LB_n      (SRAM_LB_n_from_the_sram),                         //                  .export
		.SRAM_WE_n      (SRAM_WE_n_from_the_sram),                         //                  .export
		.SRAM_CE_n      (SRAM_CE_n_from_the_sram),                         //                  .export
		.SRAM_OE_n      (SRAM_OE_n_from_the_sram)                          //                  .export
	);

	DE2_115_SOPC_sw sw (
		.clk      (altpll_0_c2_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port  (in_port_to_the_sw)                    // external_connection.export
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_0_c2_clk),                                //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_timer timer (
		.clk        (altpll_0_c2_clk),                       //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)      //   irq.irq
	);

	DE2_115_SOPC_tri_state_bridge_flash_bridge_0 tri_state_bridge_flash_bridge_0 (
		.clk                                      (altpll_0_c0_clk),                                                             //   clk.clk
		.reset                                    (rst_controller_reset_out_reset),                                              // reset.reset
		.request                                  (tri_state_bridge_flash_pinsharer_0_tcm_request),                              //   tcs.request
		.grant                                    (tri_state_bridge_flash_pinsharer_0_tcm_grant),                                //      .grant
		.tcs_data_to_and_from_the_cfi_flash       (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_out),   //      .data_to_and_from_the_cfi_flash_out
		.tcs_data_to_and_from_the_cfi_flash_outen (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_outen), //      .data_to_and_from_the_cfi_flash_outen
		.tcs_data_to_and_from_the_cfi_flash_in    (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_in),    //      .data_to_and_from_the_cfi_flash_in
		.tcs_address_to_the_cfi_flash             (tri_state_bridge_flash_pinsharer_0_tcm_address_to_the_cfi_flash_out),         //      .address_to_the_cfi_flash_out
		.tcs_write_n_to_the_cfi_flash             (tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),         //      .write_n_to_the_cfi_flash_out
		.tcs_select_n_to_the_cfi_flash            (tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),        //      .select_n_to_the_cfi_flash_out
		.tcs_read_n_to_the_cfi_flash              (tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),          //      .read_n_to_the_cfi_flash_out
		.data_to_and_from_the_cfi_flash           (data_to_and_from_the_cfi_flash),                                              //   out.data_to_and_from_the_cfi_flash
		.address_to_the_cfi_flash                 (address_to_the_cfi_flash),                                                    //      .address_to_the_cfi_flash
		.write_n_to_the_cfi_flash                 (write_n_to_the_cfi_flash),                                                    //      .write_n_to_the_cfi_flash
		.select_n_to_the_cfi_flash                (select_n_to_the_cfi_flash),                                                   //      .select_n_to_the_cfi_flash
		.read_n_to_the_cfi_flash                  (read_n_to_the_cfi_flash)                                                      //      .read_n_to_the_cfi_flash
	);

	DE2_115_SOPC_tri_state_bridge_flash_pinSharer_0 tri_state_bridge_flash_pinsharer_0 (
		.clk_clk                              (altpll_0_c0_clk),                                                             //   clk.clk
		.reset_reset                          (rst_controller_reset_out_reset),                                              // reset.reset
		.request                              (tri_state_bridge_flash_pinsharer_0_tcm_request),                              //   tcm.request
		.grant                                (tri_state_bridge_flash_pinsharer_0_tcm_grant),                                //      .grant
		.address_to_the_cfi_flash             (tri_state_bridge_flash_pinsharer_0_tcm_address_to_the_cfi_flash_out),         //      .address_to_the_cfi_flash_out
		.read_n_to_the_cfi_flash              (tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),          //      .read_n_to_the_cfi_flash_out
		.write_n_to_the_cfi_flash             (tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),         //      .write_n_to_the_cfi_flash_out
		.data_to_and_from_the_cfi_flash       (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_out),   //      .data_to_and_from_the_cfi_flash_out
		.data_to_and_from_the_cfi_flash_in    (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_in),    //      .data_to_and_from_the_cfi_flash_in
		.data_to_and_from_the_cfi_flash_outen (tri_state_bridge_flash_pinsharer_0_tcm_data_to_and_from_the_cfi_flash_outen), //      .data_to_and_from_the_cfi_flash_outen
		.select_n_to_the_cfi_flash            (tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),        //      .select_n_to_the_cfi_flash_out
		.tcs0_request                         (cfi_flash_tcm_request),                                                       //  tcs0.request
		.tcs0_grant                           (cfi_flash_tcm_grant),                                                         //      .grant
		.tcs0_address_out                     (cfi_flash_tcm_address_out),                                                   //      .address_out
		.tcs0_read_n_out                      (cfi_flash_tcm_read_n_out),                                                    //      .read_n_out
		.tcs0_write_n_out                     (cfi_flash_tcm_write_n_out),                                                   //      .write_n_out
		.tcs0_data_out                        (cfi_flash_tcm_data_out),                                                      //      .data_out
		.tcs0_data_in                         (cfi_flash_tcm_data_in),                                                       //      .data_in
		.tcs0_data_outen                      (cfi_flash_tcm_data_outen),                                                    //      .data_outen
		.tcs0_chipselect_n_out                (cfi_flash_tcm_chipselect_n_out)                                               //      .chipselect_n_out
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                                (altpll_0_c0_clk),                                                      //                                              altpll_0_c0.clk
		.altpll_0_c3_clk                                                (altpll_0_c3_clk),                                                      //                                              altpll_0_c3.clk
		.altpll_audio_c0_clk                                            (altpll_audio_c0_clk),                                                  //                                          altpll_audio_c0.clk
		.clk_50_clk_clk                                                 (clk_50),                                                               //                                               clk_50_clk.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                                       //   alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                   //     altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.altpll_audio_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                   // altpll_audio_inclk_interface_reset_reset_bridge_in_reset.reset
		.audio_clock_sink_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                                   //             audio_clock_sink_reset_reset_bridge_in_reset.reset
		.i2c_opencores_0_clock_reset_reset_bridge_in_reset_reset        (rst_controller_005_reset_out_reset),                                   //        i2c_opencores_0_clock_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                            (alt_vip_vfr_0_avalon_master_address),                                  //                              alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                        (alt_vip_vfr_0_avalon_master_waitrequest),                              //                                                         .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                         (alt_vip_vfr_0_avalon_master_burstcount),                               //                                                         .burstcount
		.alt_vip_vfr_0_avalon_master_read                               (alt_vip_vfr_0_avalon_master_read),                                     //                                                         .read
		.alt_vip_vfr_0_avalon_master_readdata                           (alt_vip_vfr_0_avalon_master_readdata),                                 //                                                         .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                      (alt_vip_vfr_0_avalon_master_readdatavalid),                            //                                                         .readdatavalid
		.cpu_data_master_address                                        (cpu_data_master_address),                                              //                                          cpu_data_master.address
		.cpu_data_master_waitrequest                                    (cpu_data_master_waitrequest),                                          //                                                         .waitrequest
		.cpu_data_master_byteenable                                     (cpu_data_master_byteenable),                                           //                                                         .byteenable
		.cpu_data_master_read                                           (cpu_data_master_read),                                                 //                                                         .read
		.cpu_data_master_readdata                                       (cpu_data_master_readdata),                                             //                                                         .readdata
		.cpu_data_master_readdatavalid                                  (cpu_data_master_readdatavalid),                                        //                                                         .readdatavalid
		.cpu_data_master_write                                          (cpu_data_master_write),                                                //                                                         .write
		.cpu_data_master_writedata                                      (cpu_data_master_writedata),                                            //                                                         .writedata
		.cpu_data_master_debugaccess                                    (cpu_data_master_debugaccess),                                          //                                                         .debugaccess
		.cpu_instruction_master_address                                 (cpu_instruction_master_address),                                       //                                   cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                             (cpu_instruction_master_waitrequest),                                   //                                                         .waitrequest
		.cpu_instruction_master_read                                    (cpu_instruction_master_read),                                          //                                                         .read
		.cpu_instruction_master_readdata                                (cpu_instruction_master_readdata),                                      //                                                         .readdata
		.cpu_instruction_master_readdatavalid                           (cpu_instruction_master_readdatavalid),                                 //                                                         .readdatavalid
		.alt_vip_vfr_0_avalon_slave_address                             (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),                 //                               alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                               (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),                   //                                                         .write
		.alt_vip_vfr_0_avalon_slave_read                                (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),                    //                                                         .read
		.alt_vip_vfr_0_avalon_slave_readdata                            (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),                //                                                         .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata),               //                                                         .writedata
		.altpll_0_pll_slave_address                                     (mm_interconnect_0_altpll_0_pll_slave_address),                         //                                       altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                       (mm_interconnect_0_altpll_0_pll_slave_write),                           //                                                         .write
		.altpll_0_pll_slave_read                                        (mm_interconnect_0_altpll_0_pll_slave_read),                            //                                                         .read
		.altpll_0_pll_slave_readdata                                    (mm_interconnect_0_altpll_0_pll_slave_readdata),                        //                                                         .readdata
		.altpll_0_pll_slave_writedata                                   (mm_interconnect_0_altpll_0_pll_slave_writedata),                       //                                                         .writedata
		.altpll_audio_pll_slave_address                                 (mm_interconnect_0_altpll_audio_pll_slave_address),                     //                                   altpll_audio_pll_slave.address
		.altpll_audio_pll_slave_write                                   (mm_interconnect_0_altpll_audio_pll_slave_write),                       //                                                         .write
		.altpll_audio_pll_slave_read                                    (mm_interconnect_0_altpll_audio_pll_slave_read),                        //                                                         .read
		.altpll_audio_pll_slave_readdata                                (mm_interconnect_0_altpll_audio_pll_slave_readdata),                    //                                                         .readdata
		.altpll_audio_pll_slave_writedata                               (mm_interconnect_0_altpll_audio_pll_slave_writedata),                   //                                                         .writedata
		.audio_avalon_slave_address                                     (mm_interconnect_0_audio_avalon_slave_address),                         //                                       audio_avalon_slave.address
		.audio_avalon_slave_write                                       (mm_interconnect_0_audio_avalon_slave_write),                           //                                                         .write
		.audio_avalon_slave_read                                        (mm_interconnect_0_audio_avalon_slave_read),                            //                                                         .read
		.audio_avalon_slave_readdata                                    (mm_interconnect_0_audio_avalon_slave_readdata),                        //                                                         .readdata
		.audio_avalon_slave_writedata                                   (mm_interconnect_0_audio_avalon_slave_writedata),                       //                                                         .writedata
		.cfi_flash_uas_address                                          (mm_interconnect_0_cfi_flash_uas_address),                              //                                            cfi_flash_uas.address
		.cfi_flash_uas_write                                            (mm_interconnect_0_cfi_flash_uas_write),                                //                                                         .write
		.cfi_flash_uas_read                                             (mm_interconnect_0_cfi_flash_uas_read),                                 //                                                         .read
		.cfi_flash_uas_readdata                                         (mm_interconnect_0_cfi_flash_uas_readdata),                             //                                                         .readdata
		.cfi_flash_uas_writedata                                        (mm_interconnect_0_cfi_flash_uas_writedata),                            //                                                         .writedata
		.cfi_flash_uas_burstcount                                       (mm_interconnect_0_cfi_flash_uas_burstcount),                           //                                                         .burstcount
		.cfi_flash_uas_byteenable                                       (mm_interconnect_0_cfi_flash_uas_byteenable),                           //                                                         .byteenable
		.cfi_flash_uas_readdatavalid                                    (mm_interconnect_0_cfi_flash_uas_readdatavalid),                        //                                                         .readdatavalid
		.cfi_flash_uas_waitrequest                                      (mm_interconnect_0_cfi_flash_uas_waitrequest),                          //                                                         .waitrequest
		.cfi_flash_uas_lock                                             (mm_interconnect_0_cfi_flash_uas_lock),                                 //                                                         .lock
		.cfi_flash_uas_debugaccess                                      (mm_interconnect_0_cfi_flash_uas_debugaccess),                          //                                                         .debugaccess
		.clock_crossing_io_s0_address                                   (mm_interconnect_0_clock_crossing_io_s0_address),                       //                                     clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                                     (mm_interconnect_0_clock_crossing_io_s0_write),                         //                                                         .write
		.clock_crossing_io_s0_read                                      (mm_interconnect_0_clock_crossing_io_s0_read),                          //                                                         .read
		.clock_crossing_io_s0_readdata                                  (mm_interconnect_0_clock_crossing_io_s0_readdata),                      //                                                         .readdata
		.clock_crossing_io_s0_writedata                                 (mm_interconnect_0_clock_crossing_io_s0_writedata),                     //                                                         .writedata
		.clock_crossing_io_s0_burstcount                                (mm_interconnect_0_clock_crossing_io_s0_burstcount),                    //                                                         .burstcount
		.clock_crossing_io_s0_byteenable                                (mm_interconnect_0_clock_crossing_io_s0_byteenable),                    //                                                         .byteenable
		.clock_crossing_io_s0_readdatavalid                             (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),                 //                                                         .readdatavalid
		.clock_crossing_io_s0_waitrequest                               (mm_interconnect_0_clock_crossing_io_s0_waitrequest),                   //                                                         .waitrequest
		.clock_crossing_io_s0_debugaccess                               (mm_interconnect_0_clock_crossing_io_s0_debugaccess),                   //                                                         .debugaccess
		.cpu_debug_mem_slave_address                                    (mm_interconnect_0_cpu_debug_mem_slave_address),                        //                                      cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                      (mm_interconnect_0_cpu_debug_mem_slave_write),                          //                                                         .write
		.cpu_debug_mem_slave_read                                       (mm_interconnect_0_cpu_debug_mem_slave_read),                           //                                                         .read
		.cpu_debug_mem_slave_readdata                                   (mm_interconnect_0_cpu_debug_mem_slave_readdata),                       //                                                         .readdata
		.cpu_debug_mem_slave_writedata                                  (mm_interconnect_0_cpu_debug_mem_slave_writedata),                      //                                                         .writedata
		.cpu_debug_mem_slave_byteenable                                 (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                     //                                                         .byteenable
		.cpu_debug_mem_slave_waitrequest                                (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                    //                                                         .waitrequest
		.cpu_debug_mem_slave_debugaccess                                (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                    //                                                         .debugaccess
		.epcs_flash_controller_epcs_control_port_address                (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    //                  epcs_flash_controller_epcs_control_port.address
		.epcs_flash_controller_epcs_control_port_write                  (mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),      //                                                         .write
		.epcs_flash_controller_epcs_control_port_read                   (mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),       //                                                         .read
		.epcs_flash_controller_epcs_control_port_readdata               (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                                                         .readdata
		.epcs_flash_controller_epcs_control_port_writedata              (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                                                         .writedata
		.epcs_flash_controller_epcs_control_port_chipselect             (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                                                         .chipselect
		.i2c_opencores_0_avalon_slave_0_address                         (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),             //                           i2c_opencores_0_avalon_slave_0.address
		.i2c_opencores_0_avalon_slave_0_write                           (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),               //                                                         .write
		.i2c_opencores_0_avalon_slave_0_readdata                        (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),            //                                                         .readdata
		.i2c_opencores_0_avalon_slave_0_writedata                       (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),           //                                                         .writedata
		.i2c_opencores_0_avalon_slave_0_waitrequest                     (~mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest),        //                                                         .waitrequest
		.i2c_opencores_0_avalon_slave_0_chipselect                      (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),          //                                                         .chipselect
		.jtag_uart_avalon_jtag_slave_address                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //                              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                                         .write
		.jtag_uart_avalon_jtag_slave_read                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                                         .read
		.jtag_uart_avalon_jtag_slave_readdata                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                                         .chipselect
		.lcd_touch_int_s1_address                                       (mm_interconnect_0_lcd_touch_int_s1_address),                           //                                         lcd_touch_int_s1.address
		.lcd_touch_int_s1_write                                         (mm_interconnect_0_lcd_touch_int_s1_write),                             //                                                         .write
		.lcd_touch_int_s1_readdata                                      (mm_interconnect_0_lcd_touch_int_s1_readdata),                          //                                                         .readdata
		.lcd_touch_int_s1_writedata                                     (mm_interconnect_0_lcd_touch_int_s1_writedata),                         //                                                         .writedata
		.lcd_touch_int_s1_chipselect                                    (mm_interconnect_0_lcd_touch_int_s1_chipselect),                        //                                                         .chipselect
		.sdram_s1_address                                               (mm_interconnect_0_sdram_s1_address),                                   //                                                 sdram_s1.address
		.sdram_s1_write                                                 (mm_interconnect_0_sdram_s1_write),                                     //                                                         .write
		.sdram_s1_read                                                  (mm_interconnect_0_sdram_s1_read),                                      //                                                         .read
		.sdram_s1_readdata                                              (mm_interconnect_0_sdram_s1_readdata),                                  //                                                         .readdata
		.sdram_s1_writedata                                             (mm_interconnect_0_sdram_s1_writedata),                                 //                                                         .writedata
		.sdram_s1_byteenable                                            (mm_interconnect_0_sdram_s1_byteenable),                                //                                                         .byteenable
		.sdram_s1_readdatavalid                                         (mm_interconnect_0_sdram_s1_readdatavalid),                             //                                                         .readdatavalid
		.sdram_s1_waitrequest                                           (mm_interconnect_0_sdram_s1_waitrequest),                               //                                                         .waitrequest
		.sdram_s1_chipselect                                            (mm_interconnect_0_sdram_s1_chipselect),                                //                                                         .chipselect
		.sram_avalon_slave_address                                      (mm_interconnect_0_sram_avalon_slave_address),                          //                                        sram_avalon_slave.address
		.sram_avalon_slave_write                                        (mm_interconnect_0_sram_avalon_slave_write),                            //                                                         .write
		.sram_avalon_slave_read                                         (mm_interconnect_0_sram_avalon_slave_read),                             //                                                         .read
		.sram_avalon_slave_readdata                                     (mm_interconnect_0_sram_avalon_slave_readdata),                         //                                                         .readdata
		.sram_avalon_slave_writedata                                    (mm_interconnect_0_sram_avalon_slave_writedata),                        //                                                         .writedata
		.sram_avalon_slave_byteenable                                   (mm_interconnect_0_sram_avalon_slave_byteenable),                       //                                                         .byteenable
		.sram_avalon_slave_chipselect                                   (mm_interconnect_0_sram_avalon_slave_chipselect)                        //                                                         .chipselect
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                                        (altpll_0_c0_clk),                                   //                                      altpll_0_c0.clk
		.altpll_0_c2_clk                                        (altpll_0_c2_clk),                                   //                                      altpll_0_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.key_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                    //                  key_reset_reset_bridge_in_reset.reset
		.sd_clk_reset_reset_bridge_in_reset_reset               (rst_controller_006_reset_out_reset),                //               sd_clk_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                      //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                  //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                   //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                   //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                         //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                     //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                        //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                    //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                  //                                                 .debugaccess
		.i2c_scl_s1_address                                     (mm_interconnect_1_i2c_scl_s1_address),              //                                       i2c_scl_s1.address
		.i2c_scl_s1_write                                       (mm_interconnect_1_i2c_scl_s1_write),                //                                                 .write
		.i2c_scl_s1_readdata                                    (mm_interconnect_1_i2c_scl_s1_readdata),             //                                                 .readdata
		.i2c_scl_s1_writedata                                   (mm_interconnect_1_i2c_scl_s1_writedata),            //                                                 .writedata
		.i2c_scl_s1_chipselect                                  (mm_interconnect_1_i2c_scl_s1_chipselect),           //                                                 .chipselect
		.i2c_sda_s1_address                                     (mm_interconnect_1_i2c_sda_s1_address),              //                                       i2c_sda_s1.address
		.i2c_sda_s1_write                                       (mm_interconnect_1_i2c_sda_s1_write),                //                                                 .write
		.i2c_sda_s1_readdata                                    (mm_interconnect_1_i2c_sda_s1_readdata),             //                                                 .readdata
		.i2c_sda_s1_writedata                                   (mm_interconnect_1_i2c_sda_s1_writedata),            //                                                 .writedata
		.i2c_sda_s1_chipselect                                  (mm_interconnect_1_i2c_sda_s1_chipselect),           //                                                 .chipselect
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),                  //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                    //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),                 //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),                //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),               //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),       //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),         //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),          //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),      //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),     //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer), //                                                 .begintransfer
		.led_s1_address                                         (mm_interconnect_1_led_s1_address),                  //                                           led_s1.address
		.led_s1_write                                           (mm_interconnect_1_led_s1_write),                    //                                                 .write
		.led_s1_readdata                                        (mm_interconnect_1_led_s1_readdata),                 //                                                 .readdata
		.led_s1_writedata                                       (mm_interconnect_1_led_s1_writedata),                //                                                 .writedata
		.led_s1_chipselect                                      (mm_interconnect_1_led_s1_chipselect),               //                                                 .chipselect
		.sd_clk_s1_address                                      (mm_interconnect_1_sd_clk_s1_address),               //                                        sd_clk_s1.address
		.sd_clk_s1_write                                        (mm_interconnect_1_sd_clk_s1_write),                 //                                                 .write
		.sd_clk_s1_readdata                                     (mm_interconnect_1_sd_clk_s1_readdata),              //                                                 .readdata
		.sd_clk_s1_writedata                                    (mm_interconnect_1_sd_clk_s1_writedata),             //                                                 .writedata
		.sd_clk_s1_chipselect                                   (mm_interconnect_1_sd_clk_s1_chipselect),            //                                                 .chipselect
		.sd_cmd_s1_address                                      (mm_interconnect_1_sd_cmd_s1_address),               //                                        sd_cmd_s1.address
		.sd_cmd_s1_write                                        (mm_interconnect_1_sd_cmd_s1_write),                 //                                                 .write
		.sd_cmd_s1_readdata                                     (mm_interconnect_1_sd_cmd_s1_readdata),              //                                                 .readdata
		.sd_cmd_s1_writedata                                    (mm_interconnect_1_sd_cmd_s1_writedata),             //                                                 .writedata
		.sd_cmd_s1_chipselect                                   (mm_interconnect_1_sd_cmd_s1_chipselect),            //                                                 .chipselect
		.sd_dat_s1_address                                      (mm_interconnect_1_sd_dat_s1_address),               //                                        sd_dat_s1.address
		.sd_dat_s1_write                                        (mm_interconnect_1_sd_dat_s1_write),                 //                                                 .write
		.sd_dat_s1_readdata                                     (mm_interconnect_1_sd_dat_s1_readdata),              //                                                 .readdata
		.sd_dat_s1_writedata                                    (mm_interconnect_1_sd_dat_s1_writedata),             //                                                 .writedata
		.sd_dat_s1_chipselect                                   (mm_interconnect_1_sd_dat_s1_chipselect),            //                                                 .chipselect
		.sd_wp_n_s1_address                                     (mm_interconnect_1_sd_wp_n_s1_address),              //                                       sd_wp_n_s1.address
		.sd_wp_n_s1_readdata                                    (mm_interconnect_1_sd_wp_n_s1_readdata),             //                                                 .readdata
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                   //                                            sw_s1.address
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),                  //                                                 .readdata
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),     //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata),    //                                                 .readdata
		.timer_s1_address                                       (mm_interconnect_1_timer_s1_address),                //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_1_timer_s1_write),                  //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_1_timer_s1_readdata),               //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_1_timer_s1_writedata),              //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_1_timer_s1_chipselect)              //                                                 .chipselect
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c3_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_005_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_0_c3_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_005_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (altpll_audio_c0_clk),                //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_0_c2_clk),                    //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (altpll_0_c3_clk),                    //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
